module tb_universal_bcd_ascii_decoder;

	wire LTR_RBO;
	wire [6:0] data;

	reg ASCII;
	reg ABI, RBI, BI, LT, AL;
	reg LC, FS, X6, X7, X9;
	reg [2:0] version;
	reg [2:0] extras;
	reg [6:0] value;

	wire D0_A, D1_D, D2_RBI, D3_BI, D4_LT, D5_C, D6_B;
	assign D0_A = ASCII ? value[0] : value[0];
	assign D1_D = ASCII ? value[1] : value[3];
	assign D2_RBI = ASCII ? value[2] : RBI;
	assign D3_BI = ASCII ? value[3] : BI;
	assign D4_LT = ASCII ? value[4] : LT;
	assign D5_C = ASCII ? value[5] : value[2];
	assign D6_B = ASCII ? value[6] : value[1];

	wire X6_x0, X9_x2, X7_x1, V0_LC, V2_ABI, V1_FS;
	assign X6_x0 = ASCII ? X6 : extras[0];
	assign X9_x2 = ASCII ? X9 : extras[2];
	assign X7_x1 = ASCII ? X7 : extras[1];
	assign V0_LC = ASCII ? LC : version[0];
	assign V2_ABI = ASCII ? ABI : version[2];
	assign V1_FS = ASCII ? FS : version[1];

	wire LTR, RBO;
	assign LTR = LTR_RBO;
	assign RBO = LTR_RBO;

	universal_bcd_ascii_decoder ubcd_ascii(
		D0_A, D1_D, D2_RBI, D3_BI, D4_LT, D5_C, D6_B,
		AL, X6_x0, X9_x2, X7_x1, V0_LC, V2_ABI, V1_FS, ASCII,
		LTR_RBO, data[4], data[3], data[2], data[1], data[0], data[6], data[5]
	);

	initial begin
		ASCII = 0;

		RBI = 1; BI = 1; LT = 1; AL = 1;

		version = 0; extras = 0;
		value = 0; #100; if (data == 7'h3F) $display("PASS 0"); else $display("FAIL 0");
		value = 1; #100; if (data == 7'h06) $display("PASS 1"); else $display("FAIL 1");
		value = 2; #100; if (data == 7'h5B) $display("PASS 2"); else $display("FAIL 2");
		value = 3; #100; if (data == 7'h4F) $display("PASS 3"); else $display("FAIL 3");
		value = 4; #100; if (data == 7'h66) $display("PASS 4"); else $display("FAIL 4");
		value = 5; #100; if (data == 7'h6D) $display("PASS 5"); else $display("FAIL 5");
		value = 6; #100; if (data == 7'h7C) $display("PASS 6"); else $display("FAIL 6");
		value = 7; #100; if (data == 7'h07) $display("PASS 7"); else $display("FAIL 7");
		value = 8; #100; if (data == 7'h7F) $display("PASS 8"); else $display("FAIL 8");
		value = 9; #100; if (data == 7'h67) $display("PASS 9"); else $display("FAIL 9");
		value = 10; #100; if (data == 7'h00) $display("PASS 10"); else $display("FAIL 10");
		value = 11; #100; if (data == 7'h00) $display("PASS 11"); else $display("FAIL 11");
		value = 12; #100; if (data == 7'h00) $display("PASS 12"); else $display("FAIL 12");
		value = 13; #100; if (data == 7'h00) $display("PASS 13"); else $display("FAIL 13");
		value = 14; #100; if (data == 7'h00) $display("PASS 14"); else $display("FAIL 14");
		value = 15; #100; if (data == 7'h00) $display("PASS 15"); else $display("FAIL 15");

		version = 1; extras = 1;
		value = 0; #100; if (data == 7'h3F) $display("PASS 0"); else $display("FAIL 0");
		value = 1; #100; if (data == 7'h06) $display("PASS 1"); else $display("FAIL 1");
		value = 2; #100; if (data == 7'h5B) $display("PASS 2"); else $display("FAIL 2");
		value = 3; #100; if (data == 7'h4F) $display("PASS 3"); else $display("FAIL 3");
		value = 4; #100; if (data == 7'h66) $display("PASS 4"); else $display("FAIL 4");
		value = 5; #100; if (data == 7'h6D) $display("PASS 5"); else $display("FAIL 5");
		value = 6; #100; if (data == 7'h7D) $display("PASS 6"); else $display("FAIL 6");
		value = 7; #100; if (data == 7'h07) $display("PASS 7"); else $display("FAIL 7");
		value = 8; #100; if (data == 7'h7F) $display("PASS 8"); else $display("FAIL 8");
		value = 9; #100; if (data == 7'h67) $display("PASS 9"); else $display("FAIL 9");
		value = 10; #100; if (data == 7'h58) $display("PASS 10"); else $display("FAIL 10");
		value = 11; #100; if (data == 7'h4C) $display("PASS 11"); else $display("FAIL 11");
		value = 12; #100; if (data == 7'h62) $display("PASS 12"); else $display("FAIL 12");
		value = 13; #100; if (data == 7'h69) $display("PASS 13"); else $display("FAIL 13");
		value = 14; #100; if (data == 7'h78) $display("PASS 14"); else $display("FAIL 14");
		value = 15; #100; if (data == 7'h00) $display("PASS 15"); else $display("FAIL 15");

		version = 2; extras = 2;
		value = 0; #100; if (data == 7'h3F) $display("PASS 0"); else $display("FAIL 0");
		value = 1; #100; if (data == 7'h06) $display("PASS 1"); else $display("FAIL 1");
		value = 2; #100; if (data == 7'h5B) $display("PASS 2"); else $display("FAIL 2");
		value = 3; #100; if (data == 7'h4F) $display("PASS 3"); else $display("FAIL 3");
		value = 4; #100; if (data == 7'h66) $display("PASS 4"); else $display("FAIL 4");
		value = 5; #100; if (data == 7'h6D) $display("PASS 5"); else $display("FAIL 5");
		value = 6; #100; if (data == 7'h7C) $display("PASS 6"); else $display("FAIL 6");
		value = 7; #100; if (data == 7'h27) $display("PASS 7"); else $display("FAIL 7");
		value = 8; #100; if (data == 7'h7F) $display("PASS 8"); else $display("FAIL 8");
		value = 9; #100; if (data == 7'h67) $display("PASS 9"); else $display("FAIL 9");
		value = 10; #100; if (data == 7'h5C) $display("PASS 10"); else $display("FAIL 10");
		value = 11; #100; if (data == 7'h63) $display("PASS 11"); else $display("FAIL 11");
		value = 12; #100; if (data == 7'h01) $display("PASS 12"); else $display("FAIL 12");
		value = 13; #100; if (data == 7'h40) $display("PASS 13"); else $display("FAIL 13");
		value = 14; #100; if (data == 7'h08) $display("PASS 14"); else $display("FAIL 14");
		value = 15; #100; if (data == 7'h00) $display("PASS 15"); else $display("FAIL 15");

		version = 3; extras = 3;
		value = 0; #100; if (data == 7'h3F) $display("PASS 0"); else $display("FAIL 0");
		value = 1; #100; if (data == 7'h06) $display("PASS 1"); else $display("FAIL 1");
		value = 2; #100; if (data == 7'h5B) $display("PASS 2"); else $display("FAIL 2");
		value = 3; #100; if (data == 7'h4F) $display("PASS 3"); else $display("FAIL 3");
		value = 4; #100; if (data == 7'h66) $display("PASS 4"); else $display("FAIL 4");
		value = 5; #100; if (data == 7'h6D) $display("PASS 5"); else $display("FAIL 5");
		value = 6; #100; if (data == 7'h7D) $display("PASS 6"); else $display("FAIL 6");
		value = 7; #100; if (data == 7'h27) $display("PASS 7"); else $display("FAIL 7");
		value = 8; #100; if (data == 7'h7F) $display("PASS 8"); else $display("FAIL 8");
		value = 9; #100; if (data == 7'h67) $display("PASS 9"); else $display("FAIL 9");
		value = 10; #100; if (data == 7'h3F) $display("PASS 10"); else $display("FAIL 10");
		value = 11; #100; if (data == 7'h06) $display("PASS 11"); else $display("FAIL 11");
		value = 12; #100; if (data == 7'h5B) $display("PASS 12"); else $display("FAIL 12");
		value = 13; #100; if (data == 7'h4F) $display("PASS 13"); else $display("FAIL 13");
		value = 14; #100; if (data == 7'h66) $display("PASS 14"); else $display("FAIL 14");
		value = 15; #100; if (data == 7'h6D) $display("PASS 15"); else $display("FAIL 15");

		version = 4; extras = 4;
		value = 0; #100; if (data == 7'h3F) $display("PASS 0"); else $display("FAIL 0");
		value = 1; #100; if (data == 7'h06) $display("PASS 1"); else $display("FAIL 1");
		value = 2; #100; if (data == 7'h5B) $display("PASS 2"); else $display("FAIL 2");
		value = 3; #100; if (data == 7'h4F) $display("PASS 3"); else $display("FAIL 3");
		value = 4; #100; if (data == 7'h66) $display("PASS 4"); else $display("FAIL 4");
		value = 5; #100; if (data == 7'h6D) $display("PASS 5"); else $display("FAIL 5");
		value = 6; #100; if (data == 7'h7C) $display("PASS 6"); else $display("FAIL 6");
		value = 7; #100; if (data == 7'h07) $display("PASS 7"); else $display("FAIL 7");
		value = 8; #100; if (data == 7'h7F) $display("PASS 8"); else $display("FAIL 8");
		value = 9; #100; if (data == 7'h6F) $display("PASS 9"); else $display("FAIL 9");
		value = 10; #100; if (data == 7'h08) $display("PASS 10"); else $display("FAIL 10");
		value = 11; #100; if (data == 7'h48) $display("PASS 11"); else $display("FAIL 11");
		value = 12; #100; if (data == 7'h49) $display("PASS 12"); else $display("FAIL 12");
		value = 13; #100; if (data == 7'h41) $display("PASS 13"); else $display("FAIL 13");
		value = 14; #100; if (data == 7'h01) $display("PASS 14"); else $display("FAIL 14");
		value = 15; #100; if (data == 7'h00) $display("PASS 15"); else $display("FAIL 15");

		version = 5; extras = 5;
		value = 0; #100; if (data == 7'h3F) $display("PASS 0"); else $display("FAIL 0");
		value = 1; #100; if (data == 7'h06) $display("PASS 1"); else $display("FAIL 1");
		value = 2; #100; if (data == 7'h5B) $display("PASS 2"); else $display("FAIL 2");
		value = 3; #100; if (data == 7'h4F) $display("PASS 3"); else $display("FAIL 3");
		value = 4; #100; if (data == 7'h66) $display("PASS 4"); else $display("FAIL 4");
		value = 5; #100; if (data == 7'h6D) $display("PASS 5"); else $display("FAIL 5");
		value = 6; #100; if (data == 7'h7D) $display("PASS 6"); else $display("FAIL 6");
		value = 7; #100; if (data == 7'h07) $display("PASS 7"); else $display("FAIL 7");
		value = 8; #100; if (data == 7'h7F) $display("PASS 8"); else $display("FAIL 8");
		value = 9; #100; if (data == 7'h6F) $display("PASS 9"); else $display("FAIL 9");
		value = 10; #100; if (data == 7'h40) $display("PASS 10"); else $display("FAIL 10");
		value = 11; #100; if (data == 7'h38) $display("PASS 11"); else $display("FAIL 11");
		value = 12; #100; if (data == 7'h39) $display("PASS 12"); else $display("FAIL 12");
		value = 13; #100; if (data == 7'h31) $display("PASS 13"); else $display("FAIL 13");
		value = 14; #100; if (data == 7'h79) $display("PASS 14"); else $display("FAIL 14");
		value = 15; #100; if (data == 7'h00) $display("PASS 15"); else $display("FAIL 15");

		version = 6; extras = 6;
		value = 0; #100; if (data == 7'h3F) $display("PASS 0"); else $display("FAIL 0");
		value = 1; #100; if (data == 7'h06) $display("PASS 1"); else $display("FAIL 1");
		value = 2; #100; if (data == 7'h5B) $display("PASS 2"); else $display("FAIL 2");
		value = 3; #100; if (data == 7'h4F) $display("PASS 3"); else $display("FAIL 3");
		value = 4; #100; if (data == 7'h66) $display("PASS 4"); else $display("FAIL 4");
		value = 5; #100; if (data == 7'h6D) $display("PASS 5"); else $display("FAIL 5");
		value = 6; #100; if (data == 7'h7C) $display("PASS 6"); else $display("FAIL 6");
		value = 7; #100; if (data == 7'h27) $display("PASS 7"); else $display("FAIL 7");
		value = 8; #100; if (data == 7'h7F) $display("PASS 8"); else $display("FAIL 8");
		value = 9; #100; if (data == 7'h6F) $display("PASS 9"); else $display("FAIL 9");
		value = 10; #100; if (data == 7'h40) $display("PASS 10"); else $display("FAIL 10");
		value = 11; #100; if (data == 7'h79) $display("PASS 11"); else $display("FAIL 11");
		value = 12; #100; if (data == 7'h76) $display("PASS 12"); else $display("FAIL 12");
		value = 13; #100; if (data == 7'h38) $display("PASS 13"); else $display("FAIL 13");
		value = 14; #100; if (data == 7'h73) $display("PASS 14"); else $display("FAIL 14");
		value = 15; #100; if (data == 7'h00) $display("PASS 15"); else $display("FAIL 15");

		version = 7; extras = 7;
		value = 0; #100; if (data == 7'h3F) $display("PASS 0"); else $display("FAIL 0");
		value = 1; #100; if (data == 7'h06) $display("PASS 1"); else $display("FAIL 1");
		value = 2; #100; if (data == 7'h5B) $display("PASS 2"); else $display("FAIL 2");
		value = 3; #100; if (data == 7'h4F) $display("PASS 3"); else $display("FAIL 3");
		value = 4; #100; if (data == 7'h66) $display("PASS 4"); else $display("FAIL 4");
		value = 5; #100; if (data == 7'h6D) $display("PASS 5"); else $display("FAIL 5");
		value = 6; #100; if (data == 7'h7D) $display("PASS 6"); else $display("FAIL 6");
		value = 7; #100; if (data == 7'h27) $display("PASS 7"); else $display("FAIL 7");
		value = 8; #100; if (data == 7'h7F) $display("PASS 8"); else $display("FAIL 8");
		value = 9; #100; if (data == 7'h6F) $display("PASS 9"); else $display("FAIL 9");
		value = 10; #100; if (data == 7'h77) $display("PASS 10"); else $display("FAIL 10");
		value = 11; #100; if (data == 7'h7C) $display("PASS 11"); else $display("FAIL 11");
		value = 12; #100; if (data == 7'h39) $display("PASS 12"); else $display("FAIL 12");
		value = 13; #100; if (data == 7'h5E) $display("PASS 13"); else $display("FAIL 13");
		value = 14; #100; if (data == 7'h79) $display("PASS 14"); else $display("FAIL 14");
		value = 15; #100; if (data == 7'h71) $display("PASS 15"); else $display("FAIL 15");

		LT = 0; #100;
		if (data == 7'h7F) $display("PASS LT"); else $display("FAIL LT");

		AL = 0; #100;
		if (data == 7'h00) $display("PASS AL"); else $display("FAIL AL");

		BI = 0; #100;
		if (data == 7'h7F) $display("PASS BI"); else $display("FAIL BI");

		ASCII = 1;

		ABI = 1; AL = 1;
		LC = 1; FS = 0;
		X6 = 1; X7 = 1; X9 = 1;

		value = 7'h20; #100; if (data == 7'h00) $display("PASS 20"); else $display("FAIL 20");
		value = 7'h21; #100; if (data == 7'h0A) $display("PASS 21"); else $display("FAIL 21");
		value = 7'h22; #100; if (data == 7'h22) $display("PASS 22"); else $display("FAIL 22");
		value = 7'h23; #100; if (data == 7'h36) $display("PASS 23"); else $display("FAIL 23");
		value = 7'h24; #100; if (data == 7'h2D) $display("PASS 24"); else $display("FAIL 24");
		value = 7'h25; #100; if (data == 7'h24) $display("PASS 25"); else $display("FAIL 25");
		value = 7'h26; #100; if (data == 7'h78) $display("PASS 26"); else $display("FAIL 26");
		value = 7'h27; #100; if (data == 7'h42) $display("PASS 27"); else $display("FAIL 27");
		value = 7'h28; #100; if (data == 7'h39) $display("PASS 28"); else $display("FAIL 28");
		value = 7'h29; #100; if (data == 7'h0F) $display("PASS 29"); else $display("FAIL 29");
		value = 7'h2A; #100; if (data == 7'h63) $display("PASS 2A"); else $display("FAIL 2A");
		value = 7'h2B; #100; if (data == 7'h46) $display("PASS 2B"); else $display("FAIL 2B");
		value = 7'h2C; #100; if (data == 7'h0C) $display("PASS 2C"); else $display("FAIL 2C");
		value = 7'h2D; #100; if (data == 7'h40) $display("PASS 2D"); else $display("FAIL 2D");
		value = 7'h2E; #100; if (data == 7'h08) $display("PASS 2E"); else $display("FAIL 2E");
		value = 7'h2F; #100; if (data == 7'h52) $display("PASS 2F"); else $display("FAIL 2F");
		value = 7'h30; #100; if (data == 7'h3F) $display("PASS 30"); else $display("FAIL 30");
		value = 7'h31; #100; if (data == 7'h06) $display("PASS 31"); else $display("FAIL 31");
		value = 7'h32; #100; if (data == 7'h5B) $display("PASS 32"); else $display("FAIL 32");
		value = 7'h33; #100; if (data == 7'h4F) $display("PASS 33"); else $display("FAIL 33");
		value = 7'h34; #100; if (data == 7'h66) $display("PASS 34"); else $display("FAIL 34");
		value = 7'h35; #100; if (data == 7'h6D) $display("PASS 35"); else $display("FAIL 35");
		value = 7'h36; #100; if (data == 7'h7D) $display("PASS 36"); else $display("FAIL 36");
		value = 7'h37; #100; if (data == 7'h27) $display("PASS 37"); else $display("FAIL 37");
		value = 7'h38; #100; if (data == 7'h7F) $display("PASS 38"); else $display("FAIL 38");
		value = 7'h39; #100; if (data == 7'h6F) $display("PASS 39"); else $display("FAIL 39");
		value = 7'h3A; #100; if (data == 7'h09) $display("PASS 3A"); else $display("FAIL 3A");
		value = 7'h3B; #100; if (data == 7'h0D) $display("PASS 3B"); else $display("FAIL 3B");
		value = 7'h3C; #100; if (data == 7'h46) $display("PASS 3C"); else $display("FAIL 3C");
		value = 7'h3D; #100; if (data == 7'h48) $display("PASS 3D"); else $display("FAIL 3D");
		value = 7'h3E; #100; if (data == 7'h70) $display("PASS 3E"); else $display("FAIL 3E");
		value = 7'h3F; #100; if (data == 7'h53) $display("PASS 3F"); else $display("FAIL 3F");
		value = 7'h40; #100; if (data == 7'h7B) $display("PASS 40"); else $display("FAIL 40");
		value = 7'h41; #100; if (data == 7'h77) $display("PASS 41"); else $display("FAIL 41");
		value = 7'h42; #100; if (data == 7'h7C) $display("PASS 42"); else $display("FAIL 42");
		value = 7'h43; #100; if (data == 7'h39) $display("PASS 43"); else $display("FAIL 43");
		value = 7'h44; #100; if (data == 7'h5E) $display("PASS 44"); else $display("FAIL 44");
		value = 7'h45; #100; if (data == 7'h79) $display("PASS 45"); else $display("FAIL 45");
		value = 7'h46; #100; if (data == 7'h71) $display("PASS 46"); else $display("FAIL 46");
		value = 7'h47; #100; if (data == 7'h3D) $display("PASS 47"); else $display("FAIL 47");
		value = 7'h48; #100; if (data == 7'h76) $display("PASS 48"); else $display("FAIL 48");
		value = 7'h49; #100; if (data == 7'h06) $display("PASS 49"); else $display("FAIL 49");
		value = 7'h4A; #100; if (data == 7'h1E) $display("PASS 4A"); else $display("FAIL 4A");
		value = 7'h4B; #100; if (data == 7'h75) $display("PASS 4B"); else $display("FAIL 4B");
		value = 7'h4C; #100; if (data == 7'h38) $display("PASS 4C"); else $display("FAIL 4C");
		value = 7'h4D; #100; if (data == 7'h2B) $display("PASS 4D"); else $display("FAIL 4D");
		value = 7'h4E; #100; if (data == 7'h37) $display("PASS 4E"); else $display("FAIL 4E");
		value = 7'h4F; #100; if (data == 7'h3F) $display("PASS 4F"); else $display("FAIL 4F");
		value = 7'h50; #100; if (data == 7'h73) $display("PASS 50"); else $display("FAIL 50");
		value = 7'h51; #100; if (data == 7'h67) $display("PASS 51"); else $display("FAIL 51");
		value = 7'h52; #100; if (data == 7'h31) $display("PASS 52"); else $display("FAIL 52");
		value = 7'h53; #100; if (data == 7'h6D) $display("PASS 53"); else $display("FAIL 53");
		value = 7'h54; #100; if (data == 7'h07) $display("PASS 54"); else $display("FAIL 54");
		value = 7'h55; #100; if (data == 7'h3E) $display("PASS 55"); else $display("FAIL 55");
		value = 7'h56; #100; if (data == 7'h6A) $display("PASS 56"); else $display("FAIL 56");
		value = 7'h57; #100; if (data == 7'h7E) $display("PASS 57"); else $display("FAIL 57");
		value = 7'h58; #100; if (data == 7'h49) $display("PASS 58"); else $display("FAIL 58");
		value = 7'h59; #100; if (data == 7'h6E) $display("PASS 59"); else $display("FAIL 59");
		value = 7'h5A; #100; if (data == 7'h5B) $display("PASS 5A"); else $display("FAIL 5A");
		value = 7'h5B; #100; if (data == 7'h39) $display("PASS 5B"); else $display("FAIL 5B");
		value = 7'h5C; #100; if (data == 7'h64) $display("PASS 5C"); else $display("FAIL 5C");
		value = 7'h5D; #100; if (data == 7'h0F) $display("PASS 5D"); else $display("FAIL 5D");
		value = 7'h5E; #100; if (data == 7'h23) $display("PASS 5E"); else $display("FAIL 5E");
		value = 7'h5F; #100; if (data == 7'h08) $display("PASS 5F"); else $display("FAIL 5F");
		value = 7'h60; #100; if (data == 7'h60) $display("PASS 60"); else $display("FAIL 60");
		value = 7'h61; #100; if (data == 7'h5F) $display("PASS 61"); else $display("FAIL 61");
		value = 7'h62; #100; if (data == 7'h7C) $display("PASS 62"); else $display("FAIL 62");
		value = 7'h63; #100; if (data == 7'h58) $display("PASS 63"); else $display("FAIL 63");
		value = 7'h64; #100; if (data == 7'h5E) $display("PASS 64"); else $display("FAIL 64");
		value = 7'h65; #100; if (data == 7'h7B) $display("PASS 65"); else $display("FAIL 65");
		value = 7'h66; #100; if (data == 7'h71) $display("PASS 66"); else $display("FAIL 66");
		value = 7'h67; #100; if (data == 7'h6F) $display("PASS 67"); else $display("FAIL 67");
		value = 7'h68; #100; if (data == 7'h74) $display("PASS 68"); else $display("FAIL 68");
		value = 7'h69; #100; if (data == 7'h05) $display("PASS 69"); else $display("FAIL 69");
		value = 7'h6A; #100; if (data == 7'h0E) $display("PASS 6A"); else $display("FAIL 6A");
		value = 7'h6B; #100; if (data == 7'h75) $display("PASS 6B"); else $display("FAIL 6B");
		value = 7'h6C; #100; if (data == 7'h06) $display("PASS 6C"); else $display("FAIL 6C");
		value = 7'h6D; #100; if (data == 7'h55) $display("PASS 6D"); else $display("FAIL 6D");
		value = 7'h6E; #100; if (data == 7'h54) $display("PASS 6E"); else $display("FAIL 6E");
		value = 7'h6F; #100; if (data == 7'h5C) $display("PASS 6F"); else $display("FAIL 6F");
		value = 7'h70; #100; if (data == 7'h73) $display("PASS 70"); else $display("FAIL 70");
		value = 7'h71; #100; if (data == 7'h67) $display("PASS 71"); else $display("FAIL 71");
		value = 7'h72; #100; if (data == 7'h50) $display("PASS 72"); else $display("FAIL 72");
		value = 7'h73; #100; if (data == 7'h6D) $display("PASS 73"); else $display("FAIL 73");
		value = 7'h74; #100; if (data == 7'h78) $display("PASS 74"); else $display("FAIL 74");
		value = 7'h75; #100; if (data == 7'h1C) $display("PASS 75"); else $display("FAIL 75");
		value = 7'h76; #100; if (data == 7'h1D) $display("PASS 76"); else $display("FAIL 76");
		value = 7'h77; #100; if (data == 7'h7E) $display("PASS 77"); else $display("FAIL 77");
		value = 7'h78; #100; if (data == 7'h48) $display("PASS 78"); else $display("FAIL 78");
		value = 7'h79; #100; if (data == 7'h6E) $display("PASS 79"); else $display("FAIL 79");
		value = 7'h7A; #100; if (data == 7'h5B) $display("PASS 7A"); else $display("FAIL 7A");
		value = 7'h7B; #100; if (data == 7'h46) $display("PASS 7B"); else $display("FAIL 7B");
		value = 7'h7C; #100; if (data == 7'h30) $display("PASS 7C"); else $display("FAIL 7C");
		value = 7'h7D; #100; if (data == 7'h70) $display("PASS 7D"); else $display("FAIL 7D");
		value = 7'h7E; #100; if (data == 7'h01) $display("PASS 7E"); else $display("FAIL 7E");
		value = 7'h7F; #100; if (data == 7'h00) $display("PASS 7F"); else $display("FAIL 7F");

		LC = 1; FS = 1;
		X6 = 0; X7 = 0; X9 = 0;

		value = 7'h20; #100; if (data == 7'h00) $display("PASS 20"); else $display("FAIL 20");
		value = 7'h21; #100; if (data == 7'h0A) $display("PASS 21"); else $display("FAIL 21");
		value = 7'h22; #100; if (data == 7'h22) $display("PASS 22"); else $display("FAIL 22");
		value = 7'h23; #100; if (data == 7'h36) $display("PASS 23"); else $display("FAIL 23");
		value = 7'h24; #100; if (data == 7'h12) $display("PASS 24"); else $display("FAIL 24");
		value = 7'h25; #100; if (data == 7'h24) $display("PASS 25"); else $display("FAIL 25");
		value = 7'h26; #100; if (data == 7'h78) $display("PASS 26"); else $display("FAIL 26");
		value = 7'h27; #100; if (data == 7'h42) $display("PASS 27"); else $display("FAIL 27");
		value = 7'h28; #100; if (data == 7'h58) $display("PASS 28"); else $display("FAIL 28");
		value = 7'h29; #100; if (data == 7'h4C) $display("PASS 29"); else $display("FAIL 29");
		value = 7'h2A; #100; if (data == 7'h63) $display("PASS 2A"); else $display("FAIL 2A");
		value = 7'h2B; #100; if (data == 7'h46) $display("PASS 2B"); else $display("FAIL 2B");
		value = 7'h2C; #100; if (data == 7'h0C) $display("PASS 2C"); else $display("FAIL 2C");
		value = 7'h2D; #100; if (data == 7'h40) $display("PASS 2D"); else $display("FAIL 2D");
		value = 7'h2E; #100; if (data == 7'h10) $display("PASS 2E"); else $display("FAIL 2E");
		value = 7'h2F; #100; if (data == 7'h52) $display("PASS 2F"); else $display("FAIL 2F");
		value = 7'h30; #100; if (data == 7'h3F) $display("PASS 30"); else $display("FAIL 30");
		value = 7'h31; #100; if (data == 7'h06) $display("PASS 31"); else $display("FAIL 31");
		value = 7'h32; #100; if (data == 7'h5B) $display("PASS 32"); else $display("FAIL 32");
		value = 7'h33; #100; if (data == 7'h4F) $display("PASS 33"); else $display("FAIL 33");
		value = 7'h34; #100; if (data == 7'h66) $display("PASS 34"); else $display("FAIL 34");
		value = 7'h35; #100; if (data == 7'h6D) $display("PASS 35"); else $display("FAIL 35");
		value = 7'h36; #100; if (data == 7'h7C) $display("PASS 36"); else $display("FAIL 36");
		value = 7'h37; #100; if (data == 7'h07) $display("PASS 37"); else $display("FAIL 37");
		value = 7'h38; #100; if (data == 7'h7F) $display("PASS 38"); else $display("FAIL 38");
		value = 7'h39; #100; if (data == 7'h67) $display("PASS 39"); else $display("FAIL 39");
		value = 7'h3A; #100; if (data == 7'h09) $display("PASS 3A"); else $display("FAIL 3A");
		value = 7'h3B; #100; if (data == 7'h0D) $display("PASS 3B"); else $display("FAIL 3B");
		value = 7'h3C; #100; if (data == 7'h61) $display("PASS 3C"); else $display("FAIL 3C");
		value = 7'h3D; #100; if (data == 7'h41) $display("PASS 3D"); else $display("FAIL 3D");
		value = 7'h3E; #100; if (data == 7'h43) $display("PASS 3E"); else $display("FAIL 3E");
		value = 7'h3F; #100; if (data == 7'h53) $display("PASS 3F"); else $display("FAIL 3F");
		value = 7'h40; #100; if (data == 7'h7B) $display("PASS 40"); else $display("FAIL 40");
		value = 7'h41; #100; if (data == 7'h77) $display("PASS 41"); else $display("FAIL 41");
		value = 7'h42; #100; if (data == 7'h7C) $display("PASS 42"); else $display("FAIL 42");
		value = 7'h43; #100; if (data == 7'h39) $display("PASS 43"); else $display("FAIL 43");
		value = 7'h44; #100; if (data == 7'h5E) $display("PASS 44"); else $display("FAIL 44");
		value = 7'h45; #100; if (data == 7'h79) $display("PASS 45"); else $display("FAIL 45");
		value = 7'h46; #100; if (data == 7'h71) $display("PASS 46"); else $display("FAIL 46");
		value = 7'h47; #100; if (data == 7'h3D) $display("PASS 47"); else $display("FAIL 47");
		value = 7'h48; #100; if (data == 7'h76) $display("PASS 48"); else $display("FAIL 48");
		value = 7'h49; #100; if (data == 7'h05) $display("PASS 49"); else $display("FAIL 49");
		value = 7'h4A; #100; if (data == 7'h1E) $display("PASS 4A"); else $display("FAIL 4A");
		value = 7'h4B; #100; if (data == 7'h75) $display("PASS 4B"); else $display("FAIL 4B");
		value = 7'h4C; #100; if (data == 7'h38) $display("PASS 4C"); else $display("FAIL 4C");
		value = 7'h4D; #100; if (data == 7'h2B) $display("PASS 4D"); else $display("FAIL 4D");
		value = 7'h4E; #100; if (data == 7'h37) $display("PASS 4E"); else $display("FAIL 4E");
		value = 7'h4F; #100; if (data == 7'h6B) $display("PASS 4F"); else $display("FAIL 4F");
		value = 7'h50; #100; if (data == 7'h73) $display("PASS 50"); else $display("FAIL 50");
		value = 7'h51; #100; if (data == 7'h67) $display("PASS 51"); else $display("FAIL 51");
		value = 7'h52; #100; if (data == 7'h31) $display("PASS 52"); else $display("FAIL 52");
		value = 7'h53; #100; if (data == 7'h2D) $display("PASS 53"); else $display("FAIL 53");
		value = 7'h54; #100; if (data == 7'h07) $display("PASS 54"); else $display("FAIL 54");
		value = 7'h55; #100; if (data == 7'h3E) $display("PASS 55"); else $display("FAIL 55");
		value = 7'h56; #100; if (data == 7'h6A) $display("PASS 56"); else $display("FAIL 56");
		value = 7'h57; #100; if (data == 7'h7E) $display("PASS 57"); else $display("FAIL 57");
		value = 7'h58; #100; if (data == 7'h49) $display("PASS 58"); else $display("FAIL 58");
		value = 7'h59; #100; if (data == 7'h6E) $display("PASS 59"); else $display("FAIL 59");
		value = 7'h5A; #100; if (data == 7'h1B) $display("PASS 5A"); else $display("FAIL 5A");
		value = 7'h5B; #100; if (data == 7'h59) $display("PASS 5B"); else $display("FAIL 5B");
		value = 7'h5C; #100; if (data == 7'h64) $display("PASS 5C"); else $display("FAIL 5C");
		value = 7'h5D; #100; if (data == 7'h4D) $display("PASS 5D"); else $display("FAIL 5D");
		value = 7'h5E; #100; if (data == 7'h23) $display("PASS 5E"); else $display("FAIL 5E");
		value = 7'h5F; #100; if (data == 7'h08) $display("PASS 5F"); else $display("FAIL 5F");
		value = 7'h60; #100; if (data == 7'h60) $display("PASS 60"); else $display("FAIL 60");
		value = 7'h61; #100; if (data == 7'h44) $display("PASS 61"); else $display("FAIL 61");
		value = 7'h62; #100; if (data == 7'h7C) $display("PASS 62"); else $display("FAIL 62");
		value = 7'h63; #100; if (data == 7'h58) $display("PASS 63"); else $display("FAIL 63");
		value = 7'h64; #100; if (data == 7'h5E) $display("PASS 64"); else $display("FAIL 64");
		value = 7'h65; #100; if (data == 7'h18) $display("PASS 65"); else $display("FAIL 65");
		value = 7'h66; #100; if (data == 7'h33) $display("PASS 66"); else $display("FAIL 66");
		value = 7'h67; #100; if (data == 7'h2F) $display("PASS 67"); else $display("FAIL 67");
		value = 7'h68; #100; if (data == 7'h74) $display("PASS 68"); else $display("FAIL 68");
		value = 7'h69; #100; if (data == 7'h05) $display("PASS 69"); else $display("FAIL 69");
		value = 7'h6A; #100; if (data == 7'h0E) $display("PASS 6A"); else $display("FAIL 6A");
		value = 7'h6B; #100; if (data == 7'h75) $display("PASS 6B"); else $display("FAIL 6B");
		value = 7'h6C; #100; if (data == 7'h3C) $display("PASS 6C"); else $display("FAIL 6C");
		value = 7'h6D; #100; if (data == 7'h55) $display("PASS 6D"); else $display("FAIL 6D");
		value = 7'h6E; #100; if (data == 7'h54) $display("PASS 6E"); else $display("FAIL 6E");
		value = 7'h6F; #100; if (data == 7'h5C) $display("PASS 6F"); else $display("FAIL 6F");
		value = 7'h70; #100; if (data == 7'h73) $display("PASS 70"); else $display("FAIL 70");
		value = 7'h71; #100; if (data == 7'h67) $display("PASS 71"); else $display("FAIL 71");
		value = 7'h72; #100; if (data == 7'h50) $display("PASS 72"); else $display("FAIL 72");
		value = 7'h73; #100; if (data == 7'h2D) $display("PASS 73"); else $display("FAIL 73");
		value = 7'h74; #100; if (data == 7'h70) $display("PASS 74"); else $display("FAIL 74");
		value = 7'h75; #100; if (data == 7'h1C) $display("PASS 75"); else $display("FAIL 75");
		value = 7'h76; #100; if (data == 7'h1D) $display("PASS 76"); else $display("FAIL 76");
		value = 7'h77; #100; if (data == 7'h7E) $display("PASS 77"); else $display("FAIL 77");
		value = 7'h78; #100; if (data == 7'h48) $display("PASS 78"); else $display("FAIL 78");
		value = 7'h79; #100; if (data == 7'h6E) $display("PASS 79"); else $display("FAIL 79");
		value = 7'h7A; #100; if (data == 7'h1B) $display("PASS 7A"); else $display("FAIL 7A");
		value = 7'h7B; #100; if (data == 7'h69) $display("PASS 7B"); else $display("FAIL 7B");
		value = 7'h7C; #100; if (data == 7'h30) $display("PASS 7C"); else $display("FAIL 7C");
		value = 7'h7D; #100; if (data == 7'h4B) $display("PASS 7D"); else $display("FAIL 7D");
		value = 7'h7E; #100; if (data == 7'h01) $display("PASS 7E"); else $display("FAIL 7E");
		value = 7'h7F; #100; if (data == 7'h00) $display("PASS 7F"); else $display("FAIL 7F");

		LC = 0; FS = 0;
		X6 = 1; X7 = 1; X9 = 1;

		value = 7'h20; #100; if (data == 7'h00) $display("PASS 20"); else $display("FAIL 20");
		value = 7'h21; #100; if (data == 7'h0A) $display("PASS 21"); else $display("FAIL 21");
		value = 7'h22; #100; if (data == 7'h22) $display("PASS 22"); else $display("FAIL 22");
		value = 7'h23; #100; if (data == 7'h36) $display("PASS 23"); else $display("FAIL 23");
		value = 7'h24; #100; if (data == 7'h2D) $display("PASS 24"); else $display("FAIL 24");
		value = 7'h25; #100; if (data == 7'h24) $display("PASS 25"); else $display("FAIL 25");
		value = 7'h26; #100; if (data == 7'h78) $display("PASS 26"); else $display("FAIL 26");
		value = 7'h27; #100; if (data == 7'h42) $display("PASS 27"); else $display("FAIL 27");
		value = 7'h28; #100; if (data == 7'h39) $display("PASS 28"); else $display("FAIL 28");
		value = 7'h29; #100; if (data == 7'h0F) $display("PASS 29"); else $display("FAIL 29");
		value = 7'h2A; #100; if (data == 7'h63) $display("PASS 2A"); else $display("FAIL 2A");
		value = 7'h2B; #100; if (data == 7'h46) $display("PASS 2B"); else $display("FAIL 2B");
		value = 7'h2C; #100; if (data == 7'h0C) $display("PASS 2C"); else $display("FAIL 2C");
		value = 7'h2D; #100; if (data == 7'h40) $display("PASS 2D"); else $display("FAIL 2D");
		value = 7'h2E; #100; if (data == 7'h08) $display("PASS 2E"); else $display("FAIL 2E");
		value = 7'h2F; #100; if (data == 7'h52) $display("PASS 2F"); else $display("FAIL 2F");
		value = 7'h30; #100; if (data == 7'h3F) $display("PASS 30"); else $display("FAIL 30");
		value = 7'h31; #100; if (data == 7'h06) $display("PASS 31"); else $display("FAIL 31");
		value = 7'h32; #100; if (data == 7'h5B) $display("PASS 32"); else $display("FAIL 32");
		value = 7'h33; #100; if (data == 7'h4F) $display("PASS 33"); else $display("FAIL 33");
		value = 7'h34; #100; if (data == 7'h66) $display("PASS 34"); else $display("FAIL 34");
		value = 7'h35; #100; if (data == 7'h6D) $display("PASS 35"); else $display("FAIL 35");
		value = 7'h36; #100; if (data == 7'h7D) $display("PASS 36"); else $display("FAIL 36");
		value = 7'h37; #100; if (data == 7'h27) $display("PASS 37"); else $display("FAIL 37");
		value = 7'h38; #100; if (data == 7'h7F) $display("PASS 38"); else $display("FAIL 38");
		value = 7'h39; #100; if (data == 7'h6F) $display("PASS 39"); else $display("FAIL 39");
		value = 7'h3A; #100; if (data == 7'h09) $display("PASS 3A"); else $display("FAIL 3A");
		value = 7'h3B; #100; if (data == 7'h0D) $display("PASS 3B"); else $display("FAIL 3B");
		value = 7'h3C; #100; if (data == 7'h46) $display("PASS 3C"); else $display("FAIL 3C");
		value = 7'h3D; #100; if (data == 7'h48) $display("PASS 3D"); else $display("FAIL 3D");
		value = 7'h3E; #100; if (data == 7'h70) $display("PASS 3E"); else $display("FAIL 3E");
		value = 7'h3F; #100; if (data == 7'h53) $display("PASS 3F"); else $display("FAIL 3F");
		value = 7'h40; #100; if (data == 7'h7B) $display("PASS 40"); else $display("FAIL 40");
		value = 7'h41; #100; if (data == 7'h77) $display("PASS 41"); else $display("FAIL 41");
		value = 7'h42; #100; if (data == 7'h7C) $display("PASS 42"); else $display("FAIL 42");
		value = 7'h43; #100; if (data == 7'h39) $display("PASS 43"); else $display("FAIL 43");
		value = 7'h44; #100; if (data == 7'h5E) $display("PASS 44"); else $display("FAIL 44");
		value = 7'h45; #100; if (data == 7'h79) $display("PASS 45"); else $display("FAIL 45");
		value = 7'h46; #100; if (data == 7'h71) $display("PASS 46"); else $display("FAIL 46");
		value = 7'h47; #100; if (data == 7'h3D) $display("PASS 47"); else $display("FAIL 47");
		value = 7'h48; #100; if (data == 7'h76) $display("PASS 48"); else $display("FAIL 48");
		value = 7'h49; #100; if (data == 7'h06) $display("PASS 49"); else $display("FAIL 49");
		value = 7'h4A; #100; if (data == 7'h1E) $display("PASS 4A"); else $display("FAIL 4A");
		value = 7'h4B; #100; if (data == 7'h75) $display("PASS 4B"); else $display("FAIL 4B");
		value = 7'h4C; #100; if (data == 7'h38) $display("PASS 4C"); else $display("FAIL 4C");
		value = 7'h4D; #100; if (data == 7'h2B) $display("PASS 4D"); else $display("FAIL 4D");
		value = 7'h4E; #100; if (data == 7'h37) $display("PASS 4E"); else $display("FAIL 4E");
		value = 7'h4F; #100; if (data == 7'h3F) $display("PASS 4F"); else $display("FAIL 4F");
		value = 7'h50; #100; if (data == 7'h73) $display("PASS 50"); else $display("FAIL 50");
		value = 7'h51; #100; if (data == 7'h67) $display("PASS 51"); else $display("FAIL 51");
		value = 7'h52; #100; if (data == 7'h31) $display("PASS 52"); else $display("FAIL 52");
		value = 7'h53; #100; if (data == 7'h6D) $display("PASS 53"); else $display("FAIL 53");
		value = 7'h54; #100; if (data == 7'h07) $display("PASS 54"); else $display("FAIL 54");
		value = 7'h55; #100; if (data == 7'h3E) $display("PASS 55"); else $display("FAIL 55");
		value = 7'h56; #100; if (data == 7'h6A) $display("PASS 56"); else $display("FAIL 56");
		value = 7'h57; #100; if (data == 7'h7E) $display("PASS 57"); else $display("FAIL 57");
		value = 7'h58; #100; if (data == 7'h49) $display("PASS 58"); else $display("FAIL 58");
		value = 7'h59; #100; if (data == 7'h6E) $display("PASS 59"); else $display("FAIL 59");
		value = 7'h5A; #100; if (data == 7'h5B) $display("PASS 5A"); else $display("FAIL 5A");
		value = 7'h5B; #100; if (data == 7'h39) $display("PASS 5B"); else $display("FAIL 5B");
		value = 7'h5C; #100; if (data == 7'h64) $display("PASS 5C"); else $display("FAIL 5C");
		value = 7'h5D; #100; if (data == 7'h0F) $display("PASS 5D"); else $display("FAIL 5D");
		value = 7'h5E; #100; if (data == 7'h23) $display("PASS 5E"); else $display("FAIL 5E");
		value = 7'h5F; #100; if (data == 7'h08) $display("PASS 5F"); else $display("FAIL 5F");
		value = 7'h60; #100; if (data == 7'h60) $display("PASS 60"); else $display("FAIL 60");
		value = 7'h61; #100; if (data == 7'h77) $display("PASS 61"); else $display("FAIL 61");
		value = 7'h62; #100; if (data == 7'h7C) $display("PASS 62"); else $display("FAIL 62");
		value = 7'h63; #100; if (data == 7'h39) $display("PASS 63"); else $display("FAIL 63");
		value = 7'h64; #100; if (data == 7'h5E) $display("PASS 64"); else $display("FAIL 64");
		value = 7'h65; #100; if (data == 7'h79) $display("PASS 65"); else $display("FAIL 65");
		value = 7'h66; #100; if (data == 7'h71) $display("PASS 66"); else $display("FAIL 66");
		value = 7'h67; #100; if (data == 7'h3D) $display("PASS 67"); else $display("FAIL 67");
		value = 7'h68; #100; if (data == 7'h76) $display("PASS 68"); else $display("FAIL 68");
		value = 7'h69; #100; if (data == 7'h06) $display("PASS 69"); else $display("FAIL 69");
		value = 7'h6A; #100; if (data == 7'h1E) $display("PASS 6A"); else $display("FAIL 6A");
		value = 7'h6B; #100; if (data == 7'h75) $display("PASS 6B"); else $display("FAIL 6B");
		value = 7'h6C; #100; if (data == 7'h38) $display("PASS 6C"); else $display("FAIL 6C");
		value = 7'h6D; #100; if (data == 7'h2B) $display("PASS 6D"); else $display("FAIL 6D");
		value = 7'h6E; #100; if (data == 7'h37) $display("PASS 6E"); else $display("FAIL 6E");
		value = 7'h6F; #100; if (data == 7'h3F) $display("PASS 6F"); else $display("FAIL 6F");
		value = 7'h70; #100; if (data == 7'h73) $display("PASS 70"); else $display("FAIL 70");
		value = 7'h71; #100; if (data == 7'h67) $display("PASS 71"); else $display("FAIL 71");
		value = 7'h72; #100; if (data == 7'h31) $display("PASS 72"); else $display("FAIL 72");
		value = 7'h73; #100; if (data == 7'h6D) $display("PASS 73"); else $display("FAIL 73");
		value = 7'h74; #100; if (data == 7'h07) $display("PASS 74"); else $display("FAIL 74");
		value = 7'h75; #100; if (data == 7'h3E) $display("PASS 75"); else $display("FAIL 75");
		value = 7'h76; #100; if (data == 7'h6A) $display("PASS 76"); else $display("FAIL 76");
		value = 7'h77; #100; if (data == 7'h7E) $display("PASS 77"); else $display("FAIL 77");
		value = 7'h78; #100; if (data == 7'h49) $display("PASS 78"); else $display("FAIL 78");
		value = 7'h79; #100; if (data == 7'h6E) $display("PASS 79"); else $display("FAIL 79");
		value = 7'h7A; #100; if (data == 7'h5B) $display("PASS 7A"); else $display("FAIL 7A");
		value = 7'h7B; #100; if (data == 7'h46) $display("PASS 7B"); else $display("FAIL 7B");
		value = 7'h7C; #100; if (data == 7'h30) $display("PASS 7C"); else $display("FAIL 7C");
		value = 7'h7D; #100; if (data == 7'h70) $display("PASS 7D"); else $display("FAIL 7D");
		value = 7'h7E; #100; if (data == 7'h01) $display("PASS 7E"); else $display("FAIL 7E");
		value = 7'h7F; #100; if (data == 7'h00) $display("PASS 7F"); else $display("FAIL 7F");

		LC = 0; FS = 1;
		X6 = 0; X7 = 0; X9 = 0;

		value = 7'h20; #100; if (data == 7'h00) $display("PASS 20"); else $display("FAIL 20");
		value = 7'h21; #100; if (data == 7'h0A) $display("PASS 21"); else $display("FAIL 21");
		value = 7'h22; #100; if (data == 7'h22) $display("PASS 22"); else $display("FAIL 22");
		value = 7'h23; #100; if (data == 7'h36) $display("PASS 23"); else $display("FAIL 23");
		value = 7'h24; #100; if (data == 7'h12) $display("PASS 24"); else $display("FAIL 24");
		value = 7'h25; #100; if (data == 7'h24) $display("PASS 25"); else $display("FAIL 25");
		value = 7'h26; #100; if (data == 7'h78) $display("PASS 26"); else $display("FAIL 26");
		value = 7'h27; #100; if (data == 7'h42) $display("PASS 27"); else $display("FAIL 27");
		value = 7'h28; #100; if (data == 7'h58) $display("PASS 28"); else $display("FAIL 28");
		value = 7'h29; #100; if (data == 7'h4C) $display("PASS 29"); else $display("FAIL 29");
		value = 7'h2A; #100; if (data == 7'h63) $display("PASS 2A"); else $display("FAIL 2A");
		value = 7'h2B; #100; if (data == 7'h46) $display("PASS 2B"); else $display("FAIL 2B");
		value = 7'h2C; #100; if (data == 7'h0C) $display("PASS 2C"); else $display("FAIL 2C");
		value = 7'h2D; #100; if (data == 7'h40) $display("PASS 2D"); else $display("FAIL 2D");
		value = 7'h2E; #100; if (data == 7'h10) $display("PASS 2E"); else $display("FAIL 2E");
		value = 7'h2F; #100; if (data == 7'h52) $display("PASS 2F"); else $display("FAIL 2F");
		value = 7'h30; #100; if (data == 7'h3F) $display("PASS 30"); else $display("FAIL 30");
		value = 7'h31; #100; if (data == 7'h06) $display("PASS 31"); else $display("FAIL 31");
		value = 7'h32; #100; if (data == 7'h5B) $display("PASS 32"); else $display("FAIL 32");
		value = 7'h33; #100; if (data == 7'h4F) $display("PASS 33"); else $display("FAIL 33");
		value = 7'h34; #100; if (data == 7'h66) $display("PASS 34"); else $display("FAIL 34");
		value = 7'h35; #100; if (data == 7'h6D) $display("PASS 35"); else $display("FAIL 35");
		value = 7'h36; #100; if (data == 7'h7C) $display("PASS 36"); else $display("FAIL 36");
		value = 7'h37; #100; if (data == 7'h07) $display("PASS 37"); else $display("FAIL 37");
		value = 7'h38; #100; if (data == 7'h7F) $display("PASS 38"); else $display("FAIL 38");
		value = 7'h39; #100; if (data == 7'h67) $display("PASS 39"); else $display("FAIL 39");
		value = 7'h3A; #100; if (data == 7'h09) $display("PASS 3A"); else $display("FAIL 3A");
		value = 7'h3B; #100; if (data == 7'h0D) $display("PASS 3B"); else $display("FAIL 3B");
		value = 7'h3C; #100; if (data == 7'h61) $display("PASS 3C"); else $display("FAIL 3C");
		value = 7'h3D; #100; if (data == 7'h41) $display("PASS 3D"); else $display("FAIL 3D");
		value = 7'h3E; #100; if (data == 7'h43) $display("PASS 3E"); else $display("FAIL 3E");
		value = 7'h3F; #100; if (data == 7'h53) $display("PASS 3F"); else $display("FAIL 3F");
		value = 7'h40; #100; if (data == 7'h7B) $display("PASS 40"); else $display("FAIL 40");
		value = 7'h41; #100; if (data == 7'h77) $display("PASS 41"); else $display("FAIL 41");
		value = 7'h42; #100; if (data == 7'h7C) $display("PASS 42"); else $display("FAIL 42");
		value = 7'h43; #100; if (data == 7'h39) $display("PASS 43"); else $display("FAIL 43");
		value = 7'h44; #100; if (data == 7'h5E) $display("PASS 44"); else $display("FAIL 44");
		value = 7'h45; #100; if (data == 7'h79) $display("PASS 45"); else $display("FAIL 45");
		value = 7'h46; #100; if (data == 7'h71) $display("PASS 46"); else $display("FAIL 46");
		value = 7'h47; #100; if (data == 7'h3D) $display("PASS 47"); else $display("FAIL 47");
		value = 7'h48; #100; if (data == 7'h76) $display("PASS 48"); else $display("FAIL 48");
		value = 7'h49; #100; if (data == 7'h05) $display("PASS 49"); else $display("FAIL 49");
		value = 7'h4A; #100; if (data == 7'h1E) $display("PASS 4A"); else $display("FAIL 4A");
		value = 7'h4B; #100; if (data == 7'h75) $display("PASS 4B"); else $display("FAIL 4B");
		value = 7'h4C; #100; if (data == 7'h38) $display("PASS 4C"); else $display("FAIL 4C");
		value = 7'h4D; #100; if (data == 7'h2B) $display("PASS 4D"); else $display("FAIL 4D");
		value = 7'h4E; #100; if (data == 7'h37) $display("PASS 4E"); else $display("FAIL 4E");
		value = 7'h4F; #100; if (data == 7'h6B) $display("PASS 4F"); else $display("FAIL 4F");
		value = 7'h50; #100; if (data == 7'h73) $display("PASS 50"); else $display("FAIL 50");
		value = 7'h51; #100; if (data == 7'h67) $display("PASS 51"); else $display("FAIL 51");
		value = 7'h52; #100; if (data == 7'h31) $display("PASS 52"); else $display("FAIL 52");
		value = 7'h53; #100; if (data == 7'h2D) $display("PASS 53"); else $display("FAIL 53");
		value = 7'h54; #100; if (data == 7'h07) $display("PASS 54"); else $display("FAIL 54");
		value = 7'h55; #100; if (data == 7'h3E) $display("PASS 55"); else $display("FAIL 55");
		value = 7'h56; #100; if (data == 7'h6A) $display("PASS 56"); else $display("FAIL 56");
		value = 7'h57; #100; if (data == 7'h7E) $display("PASS 57"); else $display("FAIL 57");
		value = 7'h58; #100; if (data == 7'h49) $display("PASS 58"); else $display("FAIL 58");
		value = 7'h59; #100; if (data == 7'h6E) $display("PASS 59"); else $display("FAIL 59");
		value = 7'h5A; #100; if (data == 7'h1B) $display("PASS 5A"); else $display("FAIL 5A");
		value = 7'h5B; #100; if (data == 7'h59) $display("PASS 5B"); else $display("FAIL 5B");
		value = 7'h5C; #100; if (data == 7'h64) $display("PASS 5C"); else $display("FAIL 5C");
		value = 7'h5D; #100; if (data == 7'h4D) $display("PASS 5D"); else $display("FAIL 5D");
		value = 7'h5E; #100; if (data == 7'h23) $display("PASS 5E"); else $display("FAIL 5E");
		value = 7'h5F; #100; if (data == 7'h08) $display("PASS 5F"); else $display("FAIL 5F");
		value = 7'h60; #100; if (data == 7'h60) $display("PASS 60"); else $display("FAIL 60");
		value = 7'h61; #100; if (data == 7'h77) $display("PASS 61"); else $display("FAIL 61");
		value = 7'h62; #100; if (data == 7'h7C) $display("PASS 62"); else $display("FAIL 62");
		value = 7'h63; #100; if (data == 7'h39) $display("PASS 63"); else $display("FAIL 63");
		value = 7'h64; #100; if (data == 7'h5E) $display("PASS 64"); else $display("FAIL 64");
		value = 7'h65; #100; if (data == 7'h79) $display("PASS 65"); else $display("FAIL 65");
		value = 7'h66; #100; if (data == 7'h71) $display("PASS 66"); else $display("FAIL 66");
		value = 7'h67; #100; if (data == 7'h3D) $display("PASS 67"); else $display("FAIL 67");
		value = 7'h68; #100; if (data == 7'h76) $display("PASS 68"); else $display("FAIL 68");
		value = 7'h69; #100; if (data == 7'h05) $display("PASS 69"); else $display("FAIL 69");
		value = 7'h6A; #100; if (data == 7'h1E) $display("PASS 6A"); else $display("FAIL 6A");
		value = 7'h6B; #100; if (data == 7'h75) $display("PASS 6B"); else $display("FAIL 6B");
		value = 7'h6C; #100; if (data == 7'h38) $display("PASS 6C"); else $display("FAIL 6C");
		value = 7'h6D; #100; if (data == 7'h2B) $display("PASS 6D"); else $display("FAIL 6D");
		value = 7'h6E; #100; if (data == 7'h37) $display("PASS 6E"); else $display("FAIL 6E");
		value = 7'h6F; #100; if (data == 7'h6B) $display("PASS 6F"); else $display("FAIL 6F");
		value = 7'h70; #100; if (data == 7'h73) $display("PASS 70"); else $display("FAIL 70");
		value = 7'h71; #100; if (data == 7'h67) $display("PASS 71"); else $display("FAIL 71");
		value = 7'h72; #100; if (data == 7'h31) $display("PASS 72"); else $display("FAIL 72");
		value = 7'h73; #100; if (data == 7'h2D) $display("PASS 73"); else $display("FAIL 73");
		value = 7'h74; #100; if (data == 7'h07) $display("PASS 74"); else $display("FAIL 74");
		value = 7'h75; #100; if (data == 7'h3E) $display("PASS 75"); else $display("FAIL 75");
		value = 7'h76; #100; if (data == 7'h6A) $display("PASS 76"); else $display("FAIL 76");
		value = 7'h77; #100; if (data == 7'h7E) $display("PASS 77"); else $display("FAIL 77");
		value = 7'h78; #100; if (data == 7'h49) $display("PASS 78"); else $display("FAIL 78");
		value = 7'h79; #100; if (data == 7'h6E) $display("PASS 79"); else $display("FAIL 79");
		value = 7'h7A; #100; if (data == 7'h1B) $display("PASS 7A"); else $display("FAIL 7A");
		value = 7'h7B; #100; if (data == 7'h69) $display("PASS 7B"); else $display("FAIL 7B");
		value = 7'h7C; #100; if (data == 7'h30) $display("PASS 7C"); else $display("FAIL 7C");
		value = 7'h7D; #100; if (data == 7'h4B) $display("PASS 7D"); else $display("FAIL 7D");
		value = 7'h7E; #100; if (data == 7'h01) $display("PASS 7E"); else $display("FAIL 7E");
		value = 7'h7F; #100; if (data == 7'h00) $display("PASS 7F"); else $display("FAIL 7F");

		ABI = 1; AL = 0; #100;
		if (data == 7'h7F) $display("PASS AL"); else $display("FAIL AL");

		ABI = 0; AL = 1; #100;
		if (data == 7'h00) $display("PASS BI"); else $display("FAIL BI");
	end

	initial begin
		$dumpfile("dump.vcd");
		$dumpvars;
	end

endmodule
