library ieee;
use ieee.std_logic_1164.all;

entity kaktovik_decoder is
	port (
		RBI, BI, LT, AL, VBI : in std_logic;
		A, B, C, D, E : in std_logic;
		RBO, V : out std_logic;
		Qa, Qb, Qc, Qd, Qe, Qf, Qg, Qh : out std_logic
	);
end entity kaktovik_decoder;

architecture kak_arch of kaktovik_decoder is
	begin
		RBO <= (A and BI) or (B and BI) or (C and BI) or (D and BI) or (E and BI) or (RBI and BI) or (BI and not LT);
		V <= (C and E) or (D and E);
		Qa <= (A and B and C and D and not AL and LT) or (A and not B and C and not D and not E and not AL and LT) or (A and not B and C and E and VBI and AL and BI) or (A and not B and not C and D and E and not AL and LT) or (A and not C and not E and AL and BI) or (not A and B and not C and D and not E and not AL and LT) or (not A and not B and C and not D and E and not AL and LT) or (not A and not B and not C and not D and not E and not AL and LT) or (not A and C and not E and AL and BI) or (not A and D and E and VBI and AL and BI) or (B and not C and E and VBI and AL and BI) or (B and not D and not E and AL and BI) or (B and not D and VBI and AL and BI) or (not B and D and not E and AL and BI) or (C and E and not VBI and not AL and LT) or (not C and not D and E and AL and BI) or (D and E and not VBI and not AL and LT) or (AL and BI and not LT) or (not AL and not BI);
		Qb <= (A and B and C and D and not AL and LT) or (A and B and not C and E and VBI and AL and BI) or (A and B and D and not E and not AL and LT) or (A and B and not D and not E and AL and BI) or (A and not B and C and not D and not AL and LT) or (A and not B and not C and D and E and not AL and LT) or (A and not C and not D and E and AL and BI) or (not A and B and C and not D and not E and not AL and LT) or (not A and B and not C and D and not AL and LT) or (not A and not B and C and not E and AL and BI) or (not A and not B and D and VBI and AL and BI) or (not A and not B and not D and E and not AL and LT) or (not A and C and D and not E and AL and BI) or (not A and C and D and VBI and AL and BI) or (B and not C and not D and AL and BI) or (B and not D and E and VBI and AL and BI) or (not B and C and D and VBI and AL and BI) or (not B and not C and not D and not E and not AL and LT) or (not B and D and not E and AL and BI) or (C and E and not VBI and not AL and LT) or (D and E and not VBI and not AL and LT) or (AL and BI and not LT) or (not AL and not BI);
		Qc <= (A and B and C and D and not AL and LT) or (A and B and not C and E and VBI and AL and BI) or (A and B and D and not E and not AL and LT) or (A and B and not D and not E and AL and BI) or (A and not B and C and not D and not AL and LT) or (A and not B and not C and D and E and not AL and LT) or (A and not B and not D and not E and not AL and LT) or (A and not C and not D and E and AL and BI) or (not A and B and C and not D and not E and not AL and LT) or (not A and B and not C and D and not AL and LT) or (not A and not B and C and not E and AL and BI) or (not A and not B and not C and not D and not RBI and not AL and LT) or (not A and not B and D and VBI and AL and BI) or (not A and not B and not D and E and not AL and LT) or (not A and not B and not E and RBI and AL and BI) or (not A and C and D and not E and AL and BI) or (not A and C and D and VBI and AL and BI) or (B and not C and not D and AL and BI) or (B and not D and E and VBI and AL and BI) or (not B and C and D and VBI and AL and BI) or (not B and D and not E and AL and BI) or (C and E and not VBI and not AL and LT) or (D and E and not VBI and not AL and LT) or (AL and BI and not LT) or (not AL and not BI);
		Qd <= (A and B and not C and not D and AL and BI) or (A and B and D and not AL and LT) or (A and B and not D and E and VBI and AL and BI) or (A and not B and C and D and VBI and AL and BI) or (A and not B and D and not E and AL and BI) or (A and C and not D and not E and not AL and LT) or (A and not C and D and E and not AL and LT) or (not A and B and C and D and not E and AL and BI) or (not A and B and C and D and VBI and AL and BI) or (not A and B and C and not D and not AL and LT) or (not A and B and not C and not E and not AL and LT) or (not A and not B and C and D and not E and not AL and LT) or (not A and not B and C and not D and not E and AL and BI) or (not A and not B and D and E and VBI and AL and BI) or (B and not C and D and not AL and LT) or (B and not C and not D and E and AL and BI) or (not B and not C and D and not E and AL and BI) or (not B and not C and not D and not AL and LT) or (not B and not D and E and not AL and LT) or (C and E and not VBI and not AL and LT) or (D and E and not VBI and not AL and LT) or (AL and BI and not LT) or (not AL and not BI);
		Qe <= (A and B and not C and not D and E and AL and BI) or (A and B and D and not AL and LT) or (A and not B and C and D and E and VBI and AL and BI) or (A and not B and not C and D and not E and AL and BI) or (A and C and not E and not AL and LT) or (A and not C and D and E and not AL and LT) or (not A and B and C and D and not E and AL and BI) or (not A and B and C and D and VBI and AL and BI) or (not A and B and not C and not AL and LT) or (not A and not B and C and D and not AL and LT) or (not A and not B and C and not D and not E and AL and BI) or (not A and not B and not C and D and E and VBI and AL and BI) or (not A and not C and not E and not AL and LT) or (B and not D and not E and not AL and LT) or (not B and not C and not D and not AL and LT) or (C and not D and E and not AL and LT) or (D and E and not VBI and not AL and LT) or (AL and BI and not LT) or (not AL and not BI);
		Qf <= (A and B and C and E and not AL and LT) or (A and not B and D and VBI and AL and BI) or (A and C and not E and AL and BI) or (not A and not B and C and not D and not AL and LT) or (not A and not B and not C and D and E and not AL and LT) or (not A and C and D and VBI and AL and BI) or (B and C and not E and AL and BI) or (B and not C and E and VBI and AL and BI) or (C and not D and E and not AL and LT) or (not C and not D and E and AL and BI) or (not C and not D and not E and not AL and LT) or (D and E and not VBI and not AL and LT) or (D and not E and AL and BI) or (AL and BI and not LT) or (not AL and not BI);
		Qg <= (A and D and E and not AL and LT) or (not A and B and C and D and VBI and AL and BI) or (not A and not B and not C and E and VBI and AL and BI) or (B and not C and D and E and not AL and LT) or (B and D and not E and AL and BI) or (not B and C and D and E and not AL and LT) or (not B and not C and not E and not AL and LT) or (C and D and not E and AL and BI) or (C and E and not VBI and not AL and LT) or (not C and not D and E and AL and BI) or (D and E and not VBI and not AL and LT) or (not D and E and VBI and AL and BI) or (not D and not E and not AL and LT) or (AL and BI and not LT) or (not AL and not BI);
		Qh <= (A and B and C and D and E and not AL and LT) or (A and B and C and D and not E and AL and BI) or (not A and E and VBI and AL and BI) or (not A and not E and not AL and LT) or (not B and E and VBI and AL and BI) or (not B and not E and not AL and LT) or (C and E and not VBI and not AL and LT) or (not C and not D and E and AL and BI) or (not C and E and VBI and AL and BI) or (not C and not E and not AL and LT) or (D and E and not VBI and not AL and LT) or (not D and E and VBI and AL and BI) or (not D and not E and not AL and LT) or (AL and BI and not LT) or (not AL and not BI);
end architecture kak_arch;
